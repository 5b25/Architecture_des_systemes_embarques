    Mac OS X            	   2   �      �                                      ATTR       �   �   *                  �     com.apple.lastuseddate#PS       �     com.dropbox.attrs    �R?a    �(    

1X��W\     �����