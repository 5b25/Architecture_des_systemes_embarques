    Mac OS X            	   2   �                                           ATTR         �   9                  �     com.apple.TextEncoding      �     com.apple.lastuseddate#PS           com.dropbox.attrs    UTF-8;134217984�R?a    �G�3    

1X��W\     �����