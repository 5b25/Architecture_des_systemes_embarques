-- DE1_SoC_QSYS.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DE1_SoC_QSYS is
	port (
		adc_ltc2308_conduit_end_CONVST   : out std_logic;                                       -- adc_ltc2308_conduit_end.CONVST
		adc_ltc2308_conduit_end_SCK      : out std_logic;                                       --                        .SCK
		adc_ltc2308_conduit_end_SDI      : out std_logic;                                       --                        .SDI
		adc_ltc2308_conduit_end_SDO      : in  std_logic                    := '0';             --                        .SDO
		avalon_pwm_inst_led_pwm_readdata : out std_logic_vector(9 downto 0);                    -- avalon_pwm_inst_led_pwm.readdata
		clk_clk                          : in  std_logic                    := '0';             --                     clk.clk
		key_external_connection_export   : in  std_logic_vector(3 downto 0) := (others => '0'); -- key_external_connection.export
		pll_sys_locked_export            : out std_logic;                                       --          pll_sys_locked.export
		pll_sys_outclk2_clk              : out std_logic;                                       --         pll_sys_outclk2.clk
		pwm_4_channel_1_qsys_writedata   : out std_logic_vector(9 downto 0);                    --    pwm_4_channel_1_qsys.writedata
		reset_reset_n                    : in  std_logic                    := '0';             --                   reset.reset_n
		seven_seg_seven_seg_pwm_hex0     : out std_logic_vector(6 downto 0);                    -- seven_seg_seven_seg_pwm.hex0
		seven_seg_seven_seg_pwm_hex1     : out std_logic_vector(6 downto 0);                    --                        .hex1
		seven_seg_seven_seg_pwm_hex2     : out std_logic_vector(6 downto 0);                    --                        .hex2
		seven_seg_seven_seg_pwm_hex3     : out std_logic_vector(6 downto 0);                    --                        .hex3
		seven_seg_seven_seg_pwm_hex4     : out std_logic_vector(6 downto 0);                    --                        .hex4
		seven_seg_seven_seg_pwm_hex5     : out std_logic_vector(6 downto 0);                    --                        .hex5
		sw_external_connection_export    : in  std_logic_vector(9 downto 0) := (others => '0')  --  sw_external_connection.export
	);
end entity DE1_SoC_QSYS;

architecture rtl of DE1_SoC_QSYS is
	component DE1_SoC_QSYS_Interval_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component DE1_SoC_QSYS_Interval_timer;

	component DE1_SoC_QSYS_KEY is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component DE1_SoC_QSYS_KEY;

	component adc_ltc2308_fifo is
		port (
			slave_chipselect_n : in  std_logic                     := 'X';             -- chipselect_n
			slave_read_n       : in  std_logic                     := 'X';             -- read_n
			slave_readdata     : out std_logic_vector(15 downto 0);                    -- readdata
			slave_addr         : in  std_logic                     := 'X';             -- address
			slave_wrtie_n      : in  std_logic                     := 'X';             -- write_n
			slave_wriredata    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			ADC_CONVST         : out std_logic;                                        -- export
			ADC_SCK            : out std_logic;                                        -- export
			ADC_SDI            : out std_logic;                                        -- export
			ADC_SDO            : in  std_logic                     := 'X';             -- export
			slave_reset_n      : in  std_logic                     := 'X';             -- reset_n
			slave_clk          : in  std_logic                     := 'X';             -- clk
			adc_clk            : in  std_logic                     := 'X'              -- clk
		);
	end component adc_ltc2308_fifo;

	component avalon_pwm is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			address    : in  std_logic                     := 'X';             -- address
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			out_port   : out std_logic_vector(9 downto 0)                      -- readdata
		);
	end component avalon_pwm;

	component DE1_SoC_QSYS_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component DE1_SoC_QSYS_jtag_uart;

	component DE1_SoC_QSYS_nios2_qsys is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(19 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(19 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component DE1_SoC_QSYS_nios2_qsys;

	component DE1_SoC_QSYS_onchip_memory2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component DE1_SoC_QSYS_onchip_memory2;

	component DE1_SoC_QSYS_pll_sys is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component DE1_SoC_QSYS_pll_sys;

	component avalon_pwm_4_channels is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			out_port   : out std_logic_vector(9 downto 0)                      -- writedata
		);
	end component avalon_pwm_4_channels;

	component DE1_SoC_sevensegs is
		port (
			clk          : in  std_logic                     := 'X';             -- clk
			reset_n      : in  std_logic                     := 'X';             -- reset_n
			address      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect_n : in  std_logic                     := 'X';             -- chipselect_n
			write_n      : in  std_logic                     := 'X';             -- write_n
			s0           : out std_logic_vector(6 downto 0);                     -- hex0
			s1           : out std_logic_vector(6 downto 0);                     -- hex1
			s2           : out std_logic_vector(6 downto 0);                     -- hex2
			s3           : out std_logic_vector(6 downto 0);                     -- hex3
			s4           : out std_logic_vector(6 downto 0);                     -- hex4
			s5           : out std_logic_vector(6 downto 0)                      -- hex5
		);
	end component DE1_SoC_sevensegs;

	component DE1_SoC_QSYS_sw is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component DE1_SoC_QSYS_sw;

	component DE1_SoC_QSYS_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component DE1_SoC_QSYS_sysid_qsys;

	component DE1_SoC_QSYS_mm_interconnect_0 is
		port (
			clk_50_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			pll_sys_outclk0_clk                               : in  std_logic                     := 'X';             -- clk
			avalon_pwm_inst_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			jtag_uart_reset_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			KEY_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			nios2_qsys_reset_n_reset_bridge_in_reset_reset    : in  std_logic                     := 'X';             -- reset
			nios2_qsys_data_master_address                    : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			nios2_qsys_data_master_waitrequest                : out std_logic;                                        -- waitrequest
			nios2_qsys_data_master_byteenable                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_qsys_data_master_read                       : in  std_logic                     := 'X';             -- read
			nios2_qsys_data_master_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_data_master_readdatavalid              : out std_logic;                                        -- readdatavalid
			nios2_qsys_data_master_write                      : in  std_logic                     := 'X';             -- write
			nios2_qsys_data_master_writedata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_data_master_debugaccess                : in  std_logic                     := 'X';             -- debugaccess
			nios2_qsys_instruction_master_address             : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			nios2_qsys_instruction_master_waitrequest         : out std_logic;                                        -- waitrequest
			nios2_qsys_instruction_master_read                : in  std_logic                     := 'X';             -- read
			nios2_qsys_instruction_master_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_instruction_master_readdatavalid       : out std_logic;                                        -- readdatavalid
			adc_ltc2308_slave_address                         : out std_logic_vector(0 downto 0);                     -- address
			adc_ltc2308_slave_write                           : out std_logic;                                        -- write
			adc_ltc2308_slave_read                            : out std_logic;                                        -- read
			adc_ltc2308_slave_readdata                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			adc_ltc2308_slave_writedata                       : out std_logic_vector(15 downto 0);                    -- writedata
			adc_ltc2308_slave_chipselect                      : out std_logic;                                        -- chipselect
			avalon_pwm_inst_avalon_slave_0_address            : out std_logic_vector(0 downto 0);                     -- address
			avalon_pwm_inst_avalon_slave_0_write              : out std_logic;                                        -- write
			avalon_pwm_inst_avalon_slave_0_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avalon_pwm_inst_avalon_slave_0_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			avalon_pwm_inst_avalon_slave_0_chipselect         : out std_logic;                                        -- chipselect
			Interval_timer_s1_address                         : out std_logic_vector(2 downto 0);                     -- address
			Interval_timer_s1_write                           : out std_logic;                                        -- write
			Interval_timer_s1_readdata                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Interval_timer_s1_writedata                       : out std_logic_vector(15 downto 0);                    -- writedata
			Interval_timer_s1_chipselect                      : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address               : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                 : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                  : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect            : out std_logic;                                        -- chipselect
			KEY_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			KEY_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_qsys_jtag_debug_module_address              : out std_logic_vector(8 downto 0);                     -- address
			nios2_qsys_jtag_debug_module_write                : out std_logic;                                        -- write
			nios2_qsys_jtag_debug_module_read                 : out std_logic;                                        -- read
			nios2_qsys_jtag_debug_module_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_qsys_jtag_debug_module_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_qsys_jtag_debug_module_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_qsys_jtag_debug_module_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			nios2_qsys_jtag_debug_module_debugaccess          : out std_logic;                                        -- debugaccess
			onchip_memory2_s1_address                         : out std_logic_vector(15 downto 0);                    -- address
			onchip_memory2_s1_write                           : out std_logic;                                        -- write
			onchip_memory2_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_s1_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_s1_chipselect                      : out std_logic;                                        -- chipselect
			onchip_memory2_s1_clken                           : out std_logic;                                        -- clken
			pwm_4_channel_1_avalon_slave_0_address            : out std_logic_vector(2 downto 0);                     -- address
			pwm_4_channel_1_avalon_slave_0_write              : out std_logic;                                        -- write
			pwm_4_channel_1_avalon_slave_0_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pwm_4_channel_1_avalon_slave_0_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			pwm_4_channel_1_avalon_slave_0_chipselect         : out std_logic;                                        -- chipselect
			seven_seg_avalon_slave_0_address                  : out std_logic_vector(3 downto 0);                     -- address
			seven_seg_avalon_slave_0_write                    : out std_logic;                                        -- write
			seven_seg_avalon_slave_0_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			seven_seg_avalon_slave_0_chipselect               : out std_logic;                                        -- chipselect
			sw_s1_address                                     : out std_logic_vector(1 downto 0);                     -- address
			sw_s1_write                                       : out std_logic;                                        -- write
			sw_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sw_s1_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			sw_s1_chipselect                                  : out std_logic;                                        -- chipselect
			sysid_qsys_control_slave_address                  : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_control_slave_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component DE1_SoC_QSYS_mm_interconnect_0;

	component DE1_SoC_QSYS_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component DE1_SoC_QSYS_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component de1_soc_qsys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component de1_soc_qsys_rst_controller;

	component de1_soc_qsys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component de1_soc_qsys_rst_controller_001;

	component de1_soc_qsys_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component de1_soc_qsys_rst_controller_002;

	component de1_soc_qsys_rst_controller_003 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component de1_soc_qsys_rst_controller_003;

	signal pll_sys_outclk0_clk                                              : std_logic;                     -- pll_sys:outclk_0 -> [adc_ltc2308:slave_clk, irq_mapper:clk, irq_synchronizer:sender_clk, jtag_uart:clk, mm_interconnect_0:pll_sys_outclk0_clk, nios2_qsys:clk, onchip_memory2:clk, rst_controller_001:clk, rst_controller_003:clk, sw:clk, sysid_qsys:clock]
	signal pll_sys_outclk1_clk                                              : std_logic;                     -- pll_sys:outclk_1 -> adc_ltc2308:adc_clk
	signal nios2_qsys_data_master_readdata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	signal nios2_qsys_data_master_waitrequest                               : std_logic;                     -- mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	signal nios2_qsys_data_master_debugaccess                               : std_logic;                     -- nios2_qsys:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	signal nios2_qsys_data_master_address                                   : std_logic_vector(19 downto 0); -- nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	signal nios2_qsys_data_master_byteenable                                : std_logic_vector(3 downto 0);  -- nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	signal nios2_qsys_data_master_read                                      : std_logic;                     -- nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	signal nios2_qsys_data_master_readdatavalid                             : std_logic;                     -- mm_interconnect_0:nios2_qsys_data_master_readdatavalid -> nios2_qsys:d_readdatavalid
	signal nios2_qsys_data_master_write                                     : std_logic;                     -- nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	signal nios2_qsys_data_master_writedata                                 : std_logic_vector(31 downto 0); -- nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	signal nios2_qsys_instruction_master_readdata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	signal nios2_qsys_instruction_master_waitrequest                        : std_logic;                     -- mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	signal nios2_qsys_instruction_master_address                            : std_logic_vector(19 downto 0); -- nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	signal nios2_qsys_instruction_master_read                               : std_logic;                     -- nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	signal nios2_qsys_instruction_master_readdatavalid                      : std_logic;                     -- mm_interconnect_0:nios2_qsys_instruction_master_readdatavalid -> nios2_qsys:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect         : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata           : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest        : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read               : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write              : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_chipselect      : std_logic;                     -- mm_interconnect_0:avalon_pwm_inst_avalon_slave_0_chipselect -> avalon_pwm_inst:chipselect
	signal mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_readdata        : std_logic_vector(31 downto 0); -- avalon_pwm_inst:readdata -> mm_interconnect_0:avalon_pwm_inst_avalon_slave_0_readdata
	signal mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:avalon_pwm_inst_avalon_slave_0_address -> avalon_pwm_inst:address
	signal mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_write           : std_logic;                     -- mm_interconnect_0:avalon_pwm_inst_avalon_slave_0_write -> mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_write:in
	signal mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:avalon_pwm_inst_avalon_slave_0_writedata -> avalon_pwm_inst:writedata
	signal mm_interconnect_0_seven_seg_avalon_slave_0_chipselect            : std_logic;                     -- mm_interconnect_0:seven_seg_avalon_slave_0_chipselect -> mm_interconnect_0_seven_seg_avalon_slave_0_chipselect:in
	signal mm_interconnect_0_seven_seg_avalon_slave_0_address               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:seven_seg_avalon_slave_0_address -> seven_seg:address
	signal mm_interconnect_0_seven_seg_avalon_slave_0_write                 : std_logic;                     -- mm_interconnect_0:seven_seg_avalon_slave_0_write -> mm_interconnect_0_seven_seg_avalon_slave_0_write:in
	signal mm_interconnect_0_seven_seg_avalon_slave_0_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:seven_seg_avalon_slave_0_writedata -> seven_seg:writedata
	signal mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_chipselect      : std_logic;                     -- mm_interconnect_0:pwm_4_channel_1_avalon_slave_0_chipselect -> pwm_4_channel_1:chipselect
	signal mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_readdata        : std_logic_vector(31 downto 0); -- pwm_4_channel_1:readdata -> mm_interconnect_0:pwm_4_channel_1_avalon_slave_0_readdata
	signal mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_address         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:pwm_4_channel_1_avalon_slave_0_address -> pwm_4_channel_1:address
	signal mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_write           : std_logic;                     -- mm_interconnect_0:pwm_4_channel_1_avalon_slave_0_write -> mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_write:in
	signal mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pwm_4_channel_1_avalon_slave_0_writedata -> pwm_4_channel_1:writedata
	signal mm_interconnect_0_sysid_qsys_control_slave_readdata              : std_logic_vector(31 downto 0); -- sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_control_slave_address               : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata          : std_logic_vector(31 downto 0); -- nios2_qsys:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_jtag_debug_module_readdata
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest       : std_logic;                     -- nios2_qsys:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_jtag_debug_module_waitrequest
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess       : std_logic;                     -- mm_interconnect_0:nios2_qsys_jtag_debug_module_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_address           : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_qsys_jtag_debug_module_address -> nios2_qsys:jtag_debug_module_address
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_read              : std_logic;                     -- mm_interconnect_0:nios2_qsys_jtag_debug_module_read -> nios2_qsys:jtag_debug_module_read
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_qsys_jtag_debug_module_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_write             : std_logic;                     -- mm_interconnect_0:nios2_qsys_jtag_debug_module_write -> nios2_qsys:jtag_debug_module_write
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_jtag_debug_module_writedata -> nios2_qsys:jtag_debug_module_writedata
	signal mm_interconnect_0_onchip_memory2_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	signal mm_interconnect_0_onchip_memory2_s1_readdata                     : std_logic_vector(31 downto 0); -- onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	signal mm_interconnect_0_onchip_memory2_s1_address                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	signal mm_interconnect_0_onchip_memory2_s1_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	signal mm_interconnect_0_onchip_memory2_s1_write                        : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	signal mm_interconnect_0_onchip_memory2_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	signal mm_interconnect_0_onchip_memory2_s1_clken                        : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	signal mm_interconnect_0_sw_s1_chipselect                               : std_logic;                     -- mm_interconnect_0:sw_s1_chipselect -> sw:chipselect
	signal mm_interconnect_0_sw_s1_readdata                                 : std_logic_vector(31 downto 0); -- sw:readdata -> mm_interconnect_0:sw_s1_readdata
	signal mm_interconnect_0_sw_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sw_s1_address -> sw:address
	signal mm_interconnect_0_sw_s1_write                                    : std_logic;                     -- mm_interconnect_0:sw_s1_write -> mm_interconnect_0_sw_s1_write:in
	signal mm_interconnect_0_sw_s1_writedata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:sw_s1_writedata -> sw:writedata
	signal mm_interconnect_0_key_s1_readdata                                : std_logic_vector(31 downto 0); -- KEY:readdata -> mm_interconnect_0:KEY_s1_readdata
	signal mm_interconnect_0_key_s1_address                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:KEY_s1_address -> KEY:address
	signal mm_interconnect_0_interval_timer_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:Interval_timer_s1_chipselect -> Interval_timer:chipselect
	signal mm_interconnect_0_interval_timer_s1_readdata                     : std_logic_vector(15 downto 0); -- Interval_timer:readdata -> mm_interconnect_0:Interval_timer_s1_readdata
	signal mm_interconnect_0_interval_timer_s1_address                      : std_logic_vector(2 downto 0);  -- mm_interconnect_0:Interval_timer_s1_address -> Interval_timer:address
	signal mm_interconnect_0_interval_timer_s1_write                        : std_logic;                     -- mm_interconnect_0:Interval_timer_s1_write -> mm_interconnect_0_interval_timer_s1_write:in
	signal mm_interconnect_0_interval_timer_s1_writedata                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:Interval_timer_s1_writedata -> Interval_timer:writedata
	signal mm_interconnect_0_adc_ltc2308_slave_chipselect                   : std_logic;                     -- mm_interconnect_0:adc_ltc2308_slave_chipselect -> mm_interconnect_0_adc_ltc2308_slave_chipselect:in
	signal mm_interconnect_0_adc_ltc2308_slave_readdata                     : std_logic_vector(15 downto 0); -- adc_ltc2308:slave_readdata -> mm_interconnect_0:adc_ltc2308_slave_readdata
	signal mm_interconnect_0_adc_ltc2308_slave_address                      : std_logic_vector(0 downto 0);  -- mm_interconnect_0:adc_ltc2308_slave_address -> adc_ltc2308:slave_addr
	signal mm_interconnect_0_adc_ltc2308_slave_read                         : std_logic;                     -- mm_interconnect_0:adc_ltc2308_slave_read -> mm_interconnect_0_adc_ltc2308_slave_read:in
	signal mm_interconnect_0_adc_ltc2308_slave_write                        : std_logic;                     -- mm_interconnect_0:adc_ltc2308_slave_write -> mm_interconnect_0_adc_ltc2308_slave_write:in
	signal mm_interconnect_0_adc_ltc2308_slave_writedata                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:adc_ltc2308_slave_writedata -> adc_ltc2308:slave_wriredata
	signal irq_mapper_receiver0_irq                                         : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                         : std_logic;                     -- sw:irq -> irq_mapper:receiver1_irq
	signal nios2_qsys_d_irq_irq                                             : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_qsys:d_irq
	signal irq_mapper_receiver2_irq                                         : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver2_irq
	signal irq_synchronizer_receiver_irq                                    : std_logic_vector(0 downto 0);  -- Interval_timer:irq -> irq_synchronizer:receiver_irq
	signal rst_controller_reset_out_reset                                   : std_logic;                     -- rst_controller:reset_out -> [irq_synchronizer:receiver_reset, mm_interconnect_0:KEY_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                               : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                           : std_logic;                     -- rst_controller_001:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	signal rst_controller_002_reset_out_reset                               : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:avalon_pwm_inst_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal nios2_qsys_jtag_debug_module_reset_reset                         : std_logic;                     -- nios2_qsys:jtag_debug_module_resetrequest -> [rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	signal rst_controller_003_reset_out_reset                               : std_logic;                     -- rst_controller_003:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:nios2_qsys_reset_n_reset_bridge_in_reset_reset, rst_controller_003_reset_out_reset:in, rst_translator_001:in_reset]
	signal rst_controller_003_reset_out_reset_req                           : std_logic;                     -- rst_controller_003:reset_req -> [nios2_qsys:reset_req, rst_translator_001:reset_req_in]
	signal reset_reset_n_ports_inv                                          : std_logic;                     -- reset_reset_n:inv -> [pll_sys:rst, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv     : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv    : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_write_ports_inv : std_logic;                     -- mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_write:inv -> avalon_pwm_inst:write_n
	signal mm_interconnect_0_seven_seg_avalon_slave_0_chipselect_ports_inv  : std_logic;                     -- mm_interconnect_0_seven_seg_avalon_slave_0_chipselect:inv -> seven_seg:chipselect_n
	signal mm_interconnect_0_seven_seg_avalon_slave_0_write_ports_inv       : std_logic;                     -- mm_interconnect_0_seven_seg_avalon_slave_0_write:inv -> seven_seg:write_n
	signal mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_write_ports_inv : std_logic;                     -- mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_write:inv -> pwm_4_channel_1:write_n
	signal mm_interconnect_0_sw_s1_write_ports_inv                          : std_logic;                     -- mm_interconnect_0_sw_s1_write:inv -> sw:write_n
	signal mm_interconnect_0_interval_timer_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_interval_timer_s1_write:inv -> Interval_timer:write_n
	signal mm_interconnect_0_adc_ltc2308_slave_chipselect_ports_inv         : std_logic;                     -- mm_interconnect_0_adc_ltc2308_slave_chipselect:inv -> adc_ltc2308:slave_chipselect_n
	signal mm_interconnect_0_adc_ltc2308_slave_read_ports_inv               : std_logic;                     -- mm_interconnect_0_adc_ltc2308_slave_read:inv -> adc_ltc2308:slave_read_n
	signal mm_interconnect_0_adc_ltc2308_slave_write_ports_inv              : std_logic;                     -- mm_interconnect_0_adc_ltc2308_slave_write:inv -> adc_ltc2308:slave_wrtie_n
	signal rst_controller_reset_out_reset_ports_inv                         : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Interval_timer:reset_n, KEY:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                     : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [adc_ltc2308:slave_reset_n, jtag_uart:rst_n, sw:reset_n, sysid_qsys:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                     : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [avalon_pwm_inst:reset_n, pwm_4_channel_1:reset_n, seven_seg:reset_n]
	signal rst_controller_003_reset_out_reset_ports_inv                     : std_logic;                     -- rst_controller_003_reset_out_reset:inv -> nios2_qsys:reset_n

begin

	interval_timer : component DE1_SoC_QSYS_Interval_timer
		port map (
			clk        => clk_clk,                                             --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            -- reset.reset_n
			address    => mm_interconnect_0_interval_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_interval_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_interval_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_interval_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_interval_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_synchronizer_receiver_irq(0)                     --   irq.irq
		);

	key : component DE1_SoC_QSYS_KEY
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_key_s1_address,         --                  s1.address
			readdata => mm_interconnect_0_key_s1_readdata,        --                    .readdata
			in_port  => key_external_connection_export            -- external_connection.export
		);

	adc_ltc2308 : component adc_ltc2308_fifo
		port map (
			slave_chipselect_n => mm_interconnect_0_adc_ltc2308_slave_chipselect_ports_inv, --          slave.chipselect_n
			slave_read_n       => mm_interconnect_0_adc_ltc2308_slave_read_ports_inv,       --               .read_n
			slave_readdata     => mm_interconnect_0_adc_ltc2308_slave_readdata,             --               .readdata
			slave_addr         => mm_interconnect_0_adc_ltc2308_slave_address(0),           --               .address
			slave_wrtie_n      => mm_interconnect_0_adc_ltc2308_slave_write_ports_inv,      --               .write_n
			slave_wriredata    => mm_interconnect_0_adc_ltc2308_slave_writedata,            --               .writedata
			ADC_CONVST         => adc_ltc2308_conduit_end_CONVST,                           --    conduit_end.export
			ADC_SCK            => adc_ltc2308_conduit_end_SCK,                              --               .export
			ADC_SDI            => adc_ltc2308_conduit_end_SDI,                              --               .export
			ADC_SDO            => adc_ltc2308_conduit_end_SDO,                              --               .export
			slave_reset_n      => rst_controller_001_reset_out_reset_ports_inv,             --     reset_sink.reset_n
			slave_clk          => pll_sys_outclk0_clk,                                      --     clock_sink.clk
			adc_clk            => pll_sys_outclk1_clk                                       -- clock_sink_adc.clk
		);

	avalon_pwm_inst : component avalon_pwm
		port map (
			clk        => clk_clk,                                                          --          clock.clk
			writedata  => mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_writedata,       -- avalon_slave_0.writedata
			chipselect => mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_chipselect,      --               .chipselect
			write_n    => mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_write_ports_inv, --               .write_n
			address    => mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_address(0),      --               .address
			readdata   => mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_readdata,        --               .readdata
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,                     --          reset.reset_n
			out_port   => avalon_pwm_inst_led_pwm_readdata                                  --        led_pwm.readdata
		);

	jtag_uart : component DE1_SoC_QSYS_jtag_uart
		port map (
			clk            => pll_sys_outclk0_clk,                                           --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	nios2_qsys : component DE1_SoC_QSYS_nios2_qsys
		port map (
			clk                                   => pll_sys_outclk0_clk,                                        --                       clk.clk
			reset_n                               => rst_controller_003_reset_out_reset_ports_inv,               --                   reset_n.reset_n
			reset_req                             => rst_controller_003_reset_out_reset_req,                     --                          .reset_req
			d_address                             => nios2_qsys_data_master_address,                             --               data_master.address
			d_byteenable                          => nios2_qsys_data_master_byteenable,                          --                          .byteenable
			d_read                                => nios2_qsys_data_master_read,                                --                          .read
			d_readdata                            => nios2_qsys_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => nios2_qsys_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => nios2_qsys_data_master_write,                               --                          .write
			d_writedata                           => nios2_qsys_data_master_writedata,                           --                          .writedata
			d_readdatavalid                       => nios2_qsys_data_master_readdatavalid,                       --                          .readdatavalid
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => nios2_qsys_instruction_master_address,                      --        instruction_master.address
			i_read                                => nios2_qsys_instruction_master_read,                         --                          .read
			i_readdata                            => nios2_qsys_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => nios2_qsys_instruction_master_waitrequest,                  --                          .waitrequest
			i_readdatavalid                       => nios2_qsys_instruction_master_readdatavalid,                --                          .readdatavalid
			d_irq                                 => nios2_qsys_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios2_qsys_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_nios2_qsys_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_nios2_qsys_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_nios2_qsys_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2 : component DE1_SoC_QSYS_onchip_memory2
		port map (
			clk        => pll_sys_outclk0_clk,                            --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req,         --       .reset_req
			freeze     => '0'                                             -- (terminated)
		);

	pll_sys : component DE1_SoC_QSYS_pll_sys
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_sys_outclk0_clk,     -- outclk0.clk
			outclk_1 => pll_sys_outclk1_clk,     -- outclk1.clk
			outclk_2 => pll_sys_outclk2_clk,     -- outclk2.clk
			locked   => pll_sys_locked_export    --  locked.export
		);

	pwm_4_channel_1 : component avalon_pwm_4_channels
		port map (
			clk        => clk_clk,                                                          --          clock.clk
			writedata  => mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_writedata,       -- avalon_slave_0.writedata
			chipselect => mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_chipselect,      --               .chipselect
			write_n    => mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_write_ports_inv, --               .write_n
			address    => mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_address,         --               .address
			readdata   => mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_readdata,        --               .readdata
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,                     --          reset.reset_n
			out_port   => pwm_4_channel_1_qsys_writedata                                    --           qsys.writedata
		);

	seven_seg : component DE1_SoC_sevensegs
		port map (
			clk          => clk_clk,                                                         --          clock.clk
			reset_n      => rst_controller_002_reset_out_reset_ports_inv,                    --          reset.reset_n
			address      => mm_interconnect_0_seven_seg_avalon_slave_0_address,              -- avalon_slave_0.address
			writedata    => mm_interconnect_0_seven_seg_avalon_slave_0_writedata,            --               .writedata
			chipselect_n => mm_interconnect_0_seven_seg_avalon_slave_0_chipselect_ports_inv, --               .chipselect_n
			write_n      => mm_interconnect_0_seven_seg_avalon_slave_0_write_ports_inv,      --               .write_n
			s0           => seven_seg_seven_seg_pwm_hex0,                                    --  seven_seg_pwm.hex0
			s1           => seven_seg_seven_seg_pwm_hex1,                                    --               .hex1
			s2           => seven_seg_seven_seg_pwm_hex2,                                    --               .hex2
			s3           => seven_seg_seven_seg_pwm_hex3,                                    --               .hex3
			s4           => seven_seg_seven_seg_pwm_hex4,                                    --               .hex4
			s5           => seven_seg_seven_seg_pwm_hex5                                     --               .hex5
		);

	sw : component DE1_SoC_QSYS_sw
		port map (
			clk        => pll_sys_outclk0_clk,                          --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_sw_s1_address,              --                  s1.address
			write_n    => mm_interconnect_0_sw_s1_write_ports_inv,      --                    .write_n
			writedata  => mm_interconnect_0_sw_s1_writedata,            --                    .writedata
			chipselect => mm_interconnect_0_sw_s1_chipselect,           --                    .chipselect
			readdata   => mm_interconnect_0_sw_s1_readdata,             --                    .readdata
			in_port    => sw_external_connection_export,                -- external_connection.export
			irq        => irq_mapper_receiver1_irq                      --                 irq.irq
		);

	sysid_qsys : component DE1_SoC_QSYS_sysid_qsys
		port map (
			clock    => pll_sys_outclk0_clk,                                   --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,          --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component DE1_SoC_QSYS_mm_interconnect_0
		port map (
			clk_50_clk_clk                                    => clk_clk,                                                     --                                  clk_50_clk.clk
			pll_sys_outclk0_clk                               => pll_sys_outclk0_clk,                                         --                             pll_sys_outclk0.clk
			avalon_pwm_inst_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                          -- avalon_pwm_inst_reset_reset_bridge_in_reset.reset
			jtag_uart_reset_reset_bridge_in_reset_reset       => rst_controller_001_reset_out_reset,                          --       jtag_uart_reset_reset_bridge_in_reset.reset
			KEY_reset_reset_bridge_in_reset_reset             => rst_controller_reset_out_reset,                              --             KEY_reset_reset_bridge_in_reset.reset
			nios2_qsys_reset_n_reset_bridge_in_reset_reset    => rst_controller_003_reset_out_reset,                          --    nios2_qsys_reset_n_reset_bridge_in_reset.reset
			nios2_qsys_data_master_address                    => nios2_qsys_data_master_address,                              --                      nios2_qsys_data_master.address
			nios2_qsys_data_master_waitrequest                => nios2_qsys_data_master_waitrequest,                          --                                            .waitrequest
			nios2_qsys_data_master_byteenable                 => nios2_qsys_data_master_byteenable,                           --                                            .byteenable
			nios2_qsys_data_master_read                       => nios2_qsys_data_master_read,                                 --                                            .read
			nios2_qsys_data_master_readdata                   => nios2_qsys_data_master_readdata,                             --                                            .readdata
			nios2_qsys_data_master_readdatavalid              => nios2_qsys_data_master_readdatavalid,                        --                                            .readdatavalid
			nios2_qsys_data_master_write                      => nios2_qsys_data_master_write,                                --                                            .write
			nios2_qsys_data_master_writedata                  => nios2_qsys_data_master_writedata,                            --                                            .writedata
			nios2_qsys_data_master_debugaccess                => nios2_qsys_data_master_debugaccess,                          --                                            .debugaccess
			nios2_qsys_instruction_master_address             => nios2_qsys_instruction_master_address,                       --               nios2_qsys_instruction_master.address
			nios2_qsys_instruction_master_waitrequest         => nios2_qsys_instruction_master_waitrequest,                   --                                            .waitrequest
			nios2_qsys_instruction_master_read                => nios2_qsys_instruction_master_read,                          --                                            .read
			nios2_qsys_instruction_master_readdata            => nios2_qsys_instruction_master_readdata,                      --                                            .readdata
			nios2_qsys_instruction_master_readdatavalid       => nios2_qsys_instruction_master_readdatavalid,                 --                                            .readdatavalid
			adc_ltc2308_slave_address                         => mm_interconnect_0_adc_ltc2308_slave_address,                 --                           adc_ltc2308_slave.address
			adc_ltc2308_slave_write                           => mm_interconnect_0_adc_ltc2308_slave_write,                   --                                            .write
			adc_ltc2308_slave_read                            => mm_interconnect_0_adc_ltc2308_slave_read,                    --                                            .read
			adc_ltc2308_slave_readdata                        => mm_interconnect_0_adc_ltc2308_slave_readdata,                --                                            .readdata
			adc_ltc2308_slave_writedata                       => mm_interconnect_0_adc_ltc2308_slave_writedata,               --                                            .writedata
			adc_ltc2308_slave_chipselect                      => mm_interconnect_0_adc_ltc2308_slave_chipselect,              --                                            .chipselect
			avalon_pwm_inst_avalon_slave_0_address            => mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_address,    --              avalon_pwm_inst_avalon_slave_0.address
			avalon_pwm_inst_avalon_slave_0_write              => mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_write,      --                                            .write
			avalon_pwm_inst_avalon_slave_0_readdata           => mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_readdata,   --                                            .readdata
			avalon_pwm_inst_avalon_slave_0_writedata          => mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_writedata,  --                                            .writedata
			avalon_pwm_inst_avalon_slave_0_chipselect         => mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_chipselect, --                                            .chipselect
			Interval_timer_s1_address                         => mm_interconnect_0_interval_timer_s1_address,                 --                           Interval_timer_s1.address
			Interval_timer_s1_write                           => mm_interconnect_0_interval_timer_s1_write,                   --                                            .write
			Interval_timer_s1_readdata                        => mm_interconnect_0_interval_timer_s1_readdata,                --                                            .readdata
			Interval_timer_s1_writedata                       => mm_interconnect_0_interval_timer_s1_writedata,               --                                            .writedata
			Interval_timer_s1_chipselect                      => mm_interconnect_0_interval_timer_s1_chipselect,              --                                            .chipselect
			jtag_uart_avalon_jtag_slave_address               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,       --                 jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,         --                                            .write
			jtag_uart_avalon_jtag_slave_read                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,          --                                            .read
			jtag_uart_avalon_jtag_slave_readdata              => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,      --                                            .readdata
			jtag_uart_avalon_jtag_slave_writedata             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,     --                                            .writedata
			jtag_uart_avalon_jtag_slave_waitrequest           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,   --                                            .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,    --                                            .chipselect
			KEY_s1_address                                    => mm_interconnect_0_key_s1_address,                            --                                      KEY_s1.address
			KEY_s1_readdata                                   => mm_interconnect_0_key_s1_readdata,                           --                                            .readdata
			nios2_qsys_jtag_debug_module_address              => mm_interconnect_0_nios2_qsys_jtag_debug_module_address,      --                nios2_qsys_jtag_debug_module.address
			nios2_qsys_jtag_debug_module_write                => mm_interconnect_0_nios2_qsys_jtag_debug_module_write,        --                                            .write
			nios2_qsys_jtag_debug_module_read                 => mm_interconnect_0_nios2_qsys_jtag_debug_module_read,         --                                            .read
			nios2_qsys_jtag_debug_module_readdata             => mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata,     --                                            .readdata
			nios2_qsys_jtag_debug_module_writedata            => mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata,    --                                            .writedata
			nios2_qsys_jtag_debug_module_byteenable           => mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable,   --                                            .byteenable
			nios2_qsys_jtag_debug_module_waitrequest          => mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest,  --                                            .waitrequest
			nios2_qsys_jtag_debug_module_debugaccess          => mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess,  --                                            .debugaccess
			onchip_memory2_s1_address                         => mm_interconnect_0_onchip_memory2_s1_address,                 --                           onchip_memory2_s1.address
			onchip_memory2_s1_write                           => mm_interconnect_0_onchip_memory2_s1_write,                   --                                            .write
			onchip_memory2_s1_readdata                        => mm_interconnect_0_onchip_memory2_s1_readdata,                --                                            .readdata
			onchip_memory2_s1_writedata                       => mm_interconnect_0_onchip_memory2_s1_writedata,               --                                            .writedata
			onchip_memory2_s1_byteenable                      => mm_interconnect_0_onchip_memory2_s1_byteenable,              --                                            .byteenable
			onchip_memory2_s1_chipselect                      => mm_interconnect_0_onchip_memory2_s1_chipselect,              --                                            .chipselect
			onchip_memory2_s1_clken                           => mm_interconnect_0_onchip_memory2_s1_clken,                   --                                            .clken
			pwm_4_channel_1_avalon_slave_0_address            => mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_address,    --              pwm_4_channel_1_avalon_slave_0.address
			pwm_4_channel_1_avalon_slave_0_write              => mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_write,      --                                            .write
			pwm_4_channel_1_avalon_slave_0_readdata           => mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_readdata,   --                                            .readdata
			pwm_4_channel_1_avalon_slave_0_writedata          => mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_writedata,  --                                            .writedata
			pwm_4_channel_1_avalon_slave_0_chipselect         => mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_chipselect, --                                            .chipselect
			seven_seg_avalon_slave_0_address                  => mm_interconnect_0_seven_seg_avalon_slave_0_address,          --                    seven_seg_avalon_slave_0.address
			seven_seg_avalon_slave_0_write                    => mm_interconnect_0_seven_seg_avalon_slave_0_write,            --                                            .write
			seven_seg_avalon_slave_0_writedata                => mm_interconnect_0_seven_seg_avalon_slave_0_writedata,        --                                            .writedata
			seven_seg_avalon_slave_0_chipselect               => mm_interconnect_0_seven_seg_avalon_slave_0_chipselect,       --                                            .chipselect
			sw_s1_address                                     => mm_interconnect_0_sw_s1_address,                             --                                       sw_s1.address
			sw_s1_write                                       => mm_interconnect_0_sw_s1_write,                               --                                            .write
			sw_s1_readdata                                    => mm_interconnect_0_sw_s1_readdata,                            --                                            .readdata
			sw_s1_writedata                                   => mm_interconnect_0_sw_s1_writedata,                           --                                            .writedata
			sw_s1_chipselect                                  => mm_interconnect_0_sw_s1_chipselect,                          --                                            .chipselect
			sysid_qsys_control_slave_address                  => mm_interconnect_0_sysid_qsys_control_slave_address,          --                    sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata                 => mm_interconnect_0_sysid_qsys_control_slave_readdata          --                                            .readdata
		);

	irq_mapper : component DE1_SoC_QSYS_irq_mapper
		port map (
			clk           => pll_sys_outclk0_clk,                --       clk.clk
			reset         => rst_controller_003_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			sender_irq    => nios2_qsys_d_irq_irq                --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_clk,                            --       receiver_clk.clk
			sender_clk     => pll_sys_outclk0_clk,                --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_003_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver2_irq            --             sender.irq
		);

	rst_controller : component de1_soc_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component de1_soc_qsys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => pll_sys_outclk0_clk,                    --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component de1_soc_qsys_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                  -- reset_in0.reset
			reset_in1      => nios2_qsys_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => clk_clk,                                  --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,       -- reset_out.reset
			reset_req      => open,                                     -- (terminated)
			reset_req_in0  => '0',                                      -- (terminated)
			reset_req_in1  => '0',                                      -- (terminated)
			reset_in2      => '0',                                      -- (terminated)
			reset_req_in2  => '0',                                      -- (terminated)
			reset_in3      => '0',                                      -- (terminated)
			reset_req_in3  => '0',                                      -- (terminated)
			reset_in4      => '0',                                      -- (terminated)
			reset_req_in4  => '0',                                      -- (terminated)
			reset_in5      => '0',                                      -- (terminated)
			reset_req_in5  => '0',                                      -- (terminated)
			reset_in6      => '0',                                      -- (terminated)
			reset_req_in6  => '0',                                      -- (terminated)
			reset_in7      => '0',                                      -- (terminated)
			reset_req_in7  => '0',                                      -- (terminated)
			reset_in8      => '0',                                      -- (terminated)
			reset_req_in8  => '0',                                      -- (terminated)
			reset_in9      => '0',                                      -- (terminated)
			reset_req_in9  => '0',                                      -- (terminated)
			reset_in10     => '0',                                      -- (terminated)
			reset_req_in10 => '0',                                      -- (terminated)
			reset_in11     => '0',                                      -- (terminated)
			reset_req_in11 => '0',                                      -- (terminated)
			reset_in12     => '0',                                      -- (terminated)
			reset_req_in12 => '0',                                      -- (terminated)
			reset_in13     => '0',                                      -- (terminated)
			reset_req_in13 => '0',                                      -- (terminated)
			reset_in14     => '0',                                      -- (terminated)
			reset_req_in14 => '0',                                      -- (terminated)
			reset_in15     => '0',                                      -- (terminated)
			reset_req_in15 => '0'                                       -- (terminated)
		);

	rst_controller_003 : component de1_soc_qsys_rst_controller_003
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                  -- reset_in0.reset
			reset_in1      => nios2_qsys_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => pll_sys_outclk0_clk,                      --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset,       -- reset_out.reset
			reset_req      => rst_controller_003_reset_out_reset_req,   --          .reset_req
			reset_req_in0  => '0',                                      -- (terminated)
			reset_req_in1  => '0',                                      -- (terminated)
			reset_in2      => '0',                                      -- (terminated)
			reset_req_in2  => '0',                                      -- (terminated)
			reset_in3      => '0',                                      -- (terminated)
			reset_req_in3  => '0',                                      -- (terminated)
			reset_in4      => '0',                                      -- (terminated)
			reset_req_in4  => '0',                                      -- (terminated)
			reset_in5      => '0',                                      -- (terminated)
			reset_req_in5  => '0',                                      -- (terminated)
			reset_in6      => '0',                                      -- (terminated)
			reset_req_in6  => '0',                                      -- (terminated)
			reset_in7      => '0',                                      -- (terminated)
			reset_req_in7  => '0',                                      -- (terminated)
			reset_in8      => '0',                                      -- (terminated)
			reset_req_in8  => '0',                                      -- (terminated)
			reset_in9      => '0',                                      -- (terminated)
			reset_req_in9  => '0',                                      -- (terminated)
			reset_in10     => '0',                                      -- (terminated)
			reset_req_in10 => '0',                                      -- (terminated)
			reset_in11     => '0',                                      -- (terminated)
			reset_req_in11 => '0',                                      -- (terminated)
			reset_in12     => '0',                                      -- (terminated)
			reset_req_in12 => '0',                                      -- (terminated)
			reset_in13     => '0',                                      -- (terminated)
			reset_req_in13 => '0',                                      -- (terminated)
			reset_in14     => '0',                                      -- (terminated)
			reset_req_in14 => '0',                                      -- (terminated)
			reset_in15     => '0',                                      -- (terminated)
			reset_req_in15 => '0'                                       -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_avalon_pwm_inst_avalon_slave_0_write;

	mm_interconnect_0_seven_seg_avalon_slave_0_chipselect_ports_inv <= not mm_interconnect_0_seven_seg_avalon_slave_0_chipselect;

	mm_interconnect_0_seven_seg_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_seven_seg_avalon_slave_0_write;

	mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_pwm_4_channel_1_avalon_slave_0_write;

	mm_interconnect_0_sw_s1_write_ports_inv <= not mm_interconnect_0_sw_s1_write;

	mm_interconnect_0_interval_timer_s1_write_ports_inv <= not mm_interconnect_0_interval_timer_s1_write;

	mm_interconnect_0_adc_ltc2308_slave_chipselect_ports_inv <= not mm_interconnect_0_adc_ltc2308_slave_chipselect;

	mm_interconnect_0_adc_ltc2308_slave_read_ports_inv <= not mm_interconnect_0_adc_ltc2308_slave_read;

	mm_interconnect_0_adc_ltc2308_slave_write_ports_inv <= not mm_interconnect_0_adc_ltc2308_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

end architecture rtl; -- of DE1_SoC_QSYS
